//AliensBusControl_TB.v
//Author: RndMnkIII. 29/12/2019. (@RndMnkIII).
//---------------------------------------------------------
//iverilog -o AliensBusControl_TB_CAPTURED_async_sim DFFasync.v PAL16L8_053326_D21.v PAL16L8_053327_D20.v AliensBusControl2.v AliensBusControl_TB_CAPTURED_async.v
//vvp AliensBusControl_TB_CAPTURED_async_sim
//gtkwave AliensBusControl_TB_CAPTURED_async.vcd
`timescale 1 ns/ 1 ps //time-unit = 1 ns, precision = 1 ps
module AliensBusControl_TB_CAPTURED_async;
    //SYSCLK=48Mhz, period 20.832ns; 12Mhz, period 83.333ns; 3Mhz period 333.33ns
	reg [16:0] x,y;

	reg AS, BK4, INIT;
	reg WOCO, RMRD;
	reg SYSCLK, NCLK12, CKE, CKQ, RWb, CRAMCS, DTAC2;
	reg [15:0] ADDR;
	wire PROG, BANK, WORK, OBJCS, VRAMCS, CRAMCSgen, IOCS, DTACgen;
	
	AliensBusControl2 ABC(.AS(AS), .BK4(BK4), .INIT(INIT), .ADRF3(ADDR[15:3]), .WOCO(WOCO), .RMRD(RMRD), .SYSCLK(SYSCLK), 
	                     .CK12_CE(~NCLK12), .NCK12_CE(NCLK12), .CKE(CKE), .CKQ(CKQ), .CKQ_CE(CKQ), .PROG(PROG), 
						 .BANK(BANK), .WORK(WORK), .OBJCS(OBJCS), .VRAMCS(VRAMCS), .CRAMCS(CRAMCSgen), .IOCS(IOCS), .DTAC(DTACgen));

	initial
	begin
		INIT=1'b1;
	end

	initial
	begin
		BK4 = 1'b0;
		RMRD = 1'b0;
		WOCO = 1'b1;
	end

	initial
	begin
		$dumpfile ("AliensBusControl_TB_CAPTURED_async.vcd");
		$dumpvars (0, AliensBusControl_TB_CAPTURED_async); //0 all variables included
		#400700 $finish;
	end
	
	
	//ADD HERE csv2testbench.py output
initial
begin
    NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; SYSCLK = 1'b1;
    #8.75; SYSCLK = 1'b0;
    #8.75; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; SYSCLK = 1'b1;
    #11.25; SYSCLK = 1'b0;
    #11.25; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; SYSCLK = 1'b1;
    #10.0; SYSCLK = 1'b0;
    #10.0; 
end
initial
begin
    CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;

end
initial
begin
    CKQ = 1'b1;
    #70.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;

end
initial
begin
    ADDR = 16'hA027;
    #230.0; ADDR = 16'hA028;
    #730.0; ADDR = 16'h9808;
    #10.0; ADDR = 16'h1A8B;
    #480.0; ADDR = 16'h228B;
    #10.0; ADDR = 16'hA029;
    #410.0; ADDR = 16'hA02A;
    #650.0; ADDR = 16'hA02E;
    #10.0; ADDR = 16'hA02F;
    #400.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA030;
    #400.0; ADDR = 16'hA031;
    #730.0; ADDR = 16'hA811;
    #10.0; ADDR = 16'h28DB;
    #320.0; ADDR = 16'h2012;
    #10.0; ADDR = 16'hA032;
    #410.0; ADDR = 16'hA033;
    #400.0; ADDR = 16'hA030;
    #10.0; ADDR = 16'hA034;
    #720.0; ADDR = 16'h9834;
    #10.0; ADDR = 16'h1A8F;
    #200.0; ADDR = 16'h1E8F;
    #10.0; ADDR = 16'h1A8F;
    #270.0; ADDR = 16'h228F;
    #10.0; ADDR = 16'hA035;
    #410.0; ADDR = 16'hA036;
    #490.0; ADDR = 16'hA037;
    #400.0; ADDR = 16'hA030;
    #10.0; ADDR = 16'hA038;
    #410.0; ADDR = 16'hA039;
    #730.0; ADDR = 16'h1A8F;
    #570.0; ADDR = 16'hA03A;
    #410.0; ADDR = 16'hA03B;
    #410.0; ADDR = 16'hA03C;
    #730.0; ADDR = 16'h1A0C;
    #10.0; ADDR = 16'h1A8D;
    #570.0; ADDR = 16'h1A8E;
    #400.0; ADDR = 16'h208E;
    #10.0; ADDR = 16'hA03D;
    #400.0; ADDR = 16'hA03C;
    #10.0; ADDR = 16'hA03E;
    #410.0; ADDR = 16'hA03F;
    #150.0; ADDR = 16'hA83F;
    #10.0; ADDR = 16'h28DB;
    #570.0; ADDR = 16'h28DC;
    #400.0; ADDR = 16'h20DC;
    #10.0; ADDR = 16'hA03F;
    #400.0; ADDR = 16'hA033;
    #10.0; ADDR = 16'hA040;
    #410.0; ADDR = 16'hA041;
    #730.0; ADDR = 16'h1A09;
    #10.0; ADDR = 16'h1A8B;
    #480.0; ADDR = 16'h1A88;
    #10.0; ADDR = 16'h1A8C;
    #110.0; ADDR = 16'h1E8C;
    #10.0; ADDR = 16'h1A8C;
    #280.0; ADDR = 16'hA042;
    #410.0; ADDR = 16'hA043;
    #490.0; ADDR = 16'hA040;
    #10.0; ADDR = 16'hA044;
    #410.0; ADDR = 16'hA045;
    #640.0; ADDR = 16'h1F45;
    #10.0; ADDR = 16'h1FED;
    #810.0; ADDR = 16'h1FEC;
    #410.0; ADDR = 16'h1FEB;
    #240.0; ADDR = 16'h27EB;
    #10.0; ADDR = 16'hA046;
    #410.0; ADDR = 16'hA047;
    #640.0; ADDR = 16'h8047;
    #10.0; ADDR = 16'h1FEC;
    #820.0; ADDR = 16'h1FED;
    #410.0; ADDR = 16'h1FEE;
    #320.0; ADDR = 16'hA04A;
    #10.0; ADDR = 16'hA048;
    #400.0; ADDR = 16'hA049;
    #410.0; ADDR = 16'hA04A;
    #160.0; ADDR = 16'h284A;
    #10.0; ADDR = 16'h28DB;
    #570.0; ADDR = 16'h28DC;
    #400.0; ADDR = 16'h20C8;
    #10.0; ADDR = 16'hA04A;
    #410.0; ADDR = 16'hA04B;
    #400.0; ADDR = 16'hA048;
    #10.0; ADDR = 16'hA04C;
    #150.0; ADDR = 16'h804C;
    #10.0; ADDR = 16'h0208;
    #740.0; ADDR = 16'h0209;
    #640.0; ADDR = 16'h0009;
    #10.0; ADDR = 16'hA04C;
    #410.0; ADDR = 16'hA04D;
    #160.0; ADDR = 16'h1FEC;
    #10.0; ADDR = 16'h1FEE;
    #400.0; ADDR = 16'h1FEF;
    #410.0; ADDR = 16'h9FD8;
    #410.0; ADDR = 16'h9FD9;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDA;
    #730.0; ADDR = 16'h1A90;
    #330.0; ADDR = 16'h9FDB;
    #410.0; ADDR = 16'h9FDC;
    #410.0; ADDR = 16'h9FDD;
    #560.0; ADDR = 16'h8FDD;
    #10.0; ADDR = 16'h08F0;
    #890.0; ADDR = 16'h08D0;
    #10.0; ADDR = 16'h9FDE;
    #410.0; ADDR = 16'h9FDF;
    #650.0; ADDR = 16'h9FD6;
    #410.0; ADDR = 16'h9FD7;
    #650.0; ADDR = 16'h1FC7;
    #10.0; ADDR = 16'h1FEF;
    #400.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h9FEE;
    #10.0; ADDR = 16'h9FEF;
    #400.0; ADDR = 16'h9FE0;
    #10.0; ADDR = 16'h9FF0;
    #400.0; ADDR = 16'h9FF1;
    #160.0; ADDR = 16'h1A90;
    #580.0; ADDR = 16'h9FF1;
    #400.0; ADDR = 16'h9FF3;
    #10.0; ADDR = 16'h9FF2;
    #240.0; ADDR = 16'h9FF3;
    #410.0; ADDR = 16'h9FF4;
    #410.0; ADDR = 16'h9FF5;
    #160.0; ADDR = 16'h1A90;
    #990.0; ADDR = 16'h9FF5;
    #400.0; ADDR = 16'h9FF6;
    #250.0; ADDR = 16'h9FF7;
    #410.0; ADDR = 16'h9FF8;
    #410.0; ADDR = 16'h9FF9;
    #730.0; ADDR = 16'h1A93;
    #490.0; ADDR = 16'h1A94;
    #410.0; ADDR = 16'h9FF8;
    #10.0; ADDR = 16'h9FFA;
    #400.0; ADDR = 16'h9FFB;
    #410.0; ADDR = 16'h9FFC;
    #730.0; ADDR = 16'h1A95;
    #500.0; ADDR = 16'h9FFD;
    #400.0; ADDR = 16'h9FFF;
    #10.0; ADDR = 16'h9FFE;
    #400.0; ADDR = 16'h9FFF;
    #740.0; ADDR = 16'h1A95;
    #490.0; ADDR = 16'hA000;
    #410.0; ADDR = 16'hA001;
    #490.0; ADDR = 16'hA000;
    #10.0; ADDR = 16'hA002;
    #400.0; ADDR = 16'hA003;
    #650.0; ADDR = 16'hA001;
    #10.0; ADDR = 16'hA015;
    #400.0; ADDR = 16'hA014;
    #10.0; ADDR = 16'hA016;
    #490.0; ADDR = 16'hA017;
    #400.0; ADDR = 16'hA010;
    #10.0; ADDR = 16'hA018;
    #410.0; ADDR = 16'hA019;
    #150.0; ADDR = 16'h9A11;
    #10.0; ADDR = 16'h1A90;
    #650.0; ADDR = 16'hA019;
    #410.0; ADDR = 16'hA01A;
    #410.0; ADDR = 16'hA01B;
    #730.0; ADDR = 16'h1A91;
    #10.0; ADDR = 16'h1A95;
    #480.0; ADDR = 16'h201C;
    #10.0; ADDR = 16'hA01C;
    #400.0; ADDR = 16'hA01D;
    #250.0; ADDR = 16'hA01E;
    #410.0; ADDR = 16'hA01F;
    #400.0; ADDR = 16'hA000;
    #10.0; ADDR = 16'hA020;
    #730.0; ADDR = 16'h2864;
    #10.0; ADDR = 16'h28E5;
    #320.0; ADDR = 16'hA021;
    #410.0; ADDR = 16'hA022;
    #410.0; ADDR = 16'hA023;
    #730.0; ADDR = 16'h2863;
    #10.0; ADDR = 16'h28E3;
    #480.0; ADDR = 16'h2020;
    #10.0; ADDR = 16'hA024;
    #410.0; ADDR = 16'hA025;
    #240.0; ADDR = 16'hA026;
    #410.0; ADDR = 16'hA027;
    #400.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA028;
    #730.0; ADDR = 16'h1A91;
    #490.0; ADDR = 16'hA029;
    #410.0; ADDR = 16'hA02A;
    #660.0; ADDR = 16'hA02F;
    #400.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA030;
    #410.0; ADDR = 16'hA031;
    #730.0; ADDR = 16'h28E1;
    #320.0; ADDR = 16'h2020;
    #10.0; ADDR = 16'hA032;
    #410.0; ADDR = 16'hA033;
    #400.0; ADDR = 16'hA030;
    #10.0; ADDR = 16'hA034;
    #720.0; ADDR = 16'h8034;
    #10.0; ADDR = 16'h1A95;
    #480.0; ADDR = 16'h1295;
    #10.0; ADDR = 16'hA035;
    #410.0; ADDR = 16'hA036;
    #490.0; ADDR = 16'hA037;
    #410.0; ADDR = 16'hA038;
    #410.0; ADDR = 16'hA039;
    #730.0; ADDR = 16'h1A15;
    #10.0; ADDR = 16'h1A95;
    #560.0; ADDR = 16'h2090;
    #10.0; ADDR = 16'hA03A;
    #400.0; ADDR = 16'hA03B;
    #410.0; ADDR = 16'hA038;
    #10.0; ADDR = 16'hA03C;
    #720.0; ADDR = 16'h803C;
    #10.0; ADDR = 16'h1A93;
    #570.0; ADDR = 16'h1A94;
    #410.0; ADDR = 16'hA03D;
    #410.0; ADDR = 16'hA03E;
    #410.0; ADDR = 16'hA03F;
    #160.0; ADDR = 16'h28E1;
    #570.0; ADDR = 16'h28E0;
    #10.0; ADDR = 16'h28E2;
    #400.0; ADDR = 16'hA03F;
    #410.0; ADDR = 16'hA000;
    #10.0; ADDR = 16'hA040;
    #400.0; ADDR = 16'hA041;
    #730.0; ADDR = 16'h1A01;
    #10.0; ADDR = 16'h1A91;
    #490.0; ADDR = 16'h1A92;
    #400.0; ADDR = 16'h2042;
    #10.0; ADDR = 16'hA042;
    #400.0; ADDR = 16'hA043;
    #490.0; ADDR = 16'hA040;
    #10.0; ADDR = 16'hA044;
    #410.0; ADDR = 16'hA045;
    #640.0; ADDR = 16'h9845;
    #10.0; ADDR = 16'h1FED;
    #810.0; ADDR = 16'h1FEC;
    #410.0; ADDR = 16'h1FE8;
    #10.0; ADDR = 16'h1FEB;
    #240.0; ADDR = 16'hA046;
    #410.0; ADDR = 16'hA047;
    #650.0; ADDR = 16'h1F4C;
    #10.0; ADDR = 16'h1FEC;
    #810.0; ADDR = 16'h1FED;
    #410.0; ADDR = 16'h1FEE;
    #320.0; ADDR = 16'h20EE;
    #10.0; ADDR = 16'hA048;
    #410.0; ADDR = 16'hA049;
    #400.0; ADDR = 16'hA048;
    #10.0; ADDR = 16'hA04A;
    #160.0; ADDR = 16'h28E1;
    #570.0; ADDR = 16'h28E2;
    #400.0; ADDR = 16'h20E2;
    #10.0; ADDR = 16'hA04A;
    #410.0; ADDR = 16'hA04B;
    #400.0; ADDR = 16'hA049;
    #10.0; ADDR = 16'hA04C;
    #160.0; ADDR = 16'h020A;
    #900.0; ADDR = 16'h020B;
    #650.0; ADDR = 16'h2008;
    #10.0; ADDR = 16'hA04C;
    #410.0; ADDR = 16'hA04D;
    #150.0; ADDR = 16'h804D;
    #10.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h1FEF;
    #400.0; ADDR = 16'h1FE8;
    #10.0; ADDR = 16'h9FD8;
    #410.0; ADDR = 16'h9FD9;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDA;
    #730.0; ADDR = 16'h1A96;
    #320.0; ADDR = 16'h1A92;
    #10.0; ADDR = 16'h9FDB;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDC;
    #410.0; ADDR = 16'h9FDD;
    #560.0; ADDR = 16'h8FFD;
    #10.0; ADDR = 16'h08F0;
    #890.0; ADDR = 16'h08D0;
    #10.0; ADDR = 16'h9FDE;
    #400.0; ADDR = 16'h9FDF;
    #660.0; ADDR = 16'h9FD6;
    #410.0; ADDR = 16'h9FD7;
    #650.0; ADDR = 16'h1FEF;
    #410.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h9FEF;
    #410.0; ADDR = 16'h9FF0;
    #410.0; ADDR = 16'h9FF1;
    #160.0; ADDR = 16'h1A96;
    #570.0; ADDR = 16'h1B90;
    #10.0; ADDR = 16'h9FF1;
    #400.0; ADDR = 16'h9FF2;
    #250.0; ADDR = 16'h9FF3;
    #410.0; ADDR = 16'h9FF4;
    #410.0; ADDR = 16'h9FF5;
    #160.0; ADDR = 16'h1A96;
    #980.0; ADDR = 16'h9FF4;
    #10.0; ADDR = 16'h9FF5;
    #400.0; ADDR = 16'h9FF6;
    #250.0; ADDR = 16'h9FF7;
    #400.0; ADDR = 16'h9FF8;
    #420.0; ADDR = 16'h9FF9;
    #730.0; ADDR = 16'h1A99;
    #490.0; ADDR = 16'h1A9A;
    #410.0; ADDR = 16'h9FFA;
    #410.0; ADDR = 16'h9FFB;
    #400.0; ADDR = 16'h9FF8;
    #10.0; ADDR = 16'h9FFC;
    #730.0; ADDR = 16'h1A9B;
    #490.0; ADDR = 16'h9FFD;
    #410.0; ADDR = 16'h9FFE;
    #410.0; ADDR = 16'h9FFF;
    #730.0; ADDR = 16'h1A9B;
    #490.0; ADDR = 16'h2083;
    #10.0; ADDR = 16'hA000;
    #400.0; ADDR = 16'hA001;
    #490.0; ADDR = 16'hA000;
    #10.0; ADDR = 16'hA002;
    #410.0; ADDR = 16'hA003;
    #650.0; ADDR = 16'hA015;
    #400.0; ADDR = 16'hA014;
    #10.0; ADDR = 16'hA016;
    #490.0; ADDR = 16'hA017;
    #400.0; ADDR = 16'hA010;
    #10.0; ADDR = 16'hA018;
    #410.0; ADDR = 16'hA019;
    #150.0; ADDR = 16'h9819;
    #10.0; ADDR = 16'h1A96;
    #650.0; ADDR = 16'hA019;
    #410.0; ADDR = 16'hA01A;
    #410.0; ADDR = 16'hA01B;
    #730.0; ADDR = 16'h9A1B;
    #10.0; ADDR = 16'h1A9B;
    #480.0; ADDR = 16'h209B;
    #10.0; ADDR = 16'hA01C;
    #400.0; ADDR = 16'hA01D;
    #250.0; ADDR = 16'hA01C;
    #10.0; ADDR = 16'hA01E;
    #400.0; ADDR = 16'hA01F;
    #410.0; ADDR = 16'hA020;
    #730.0; ADDR = 16'hA820;
    #10.0; ADDR = 16'h28EB;
    #320.0; ADDR = 16'hA021;
    #410.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA022;
    #400.0; ADDR = 16'hA023;
    #730.0; ADDR = 16'hA823;
    #10.0; ADDR = 16'h28E9;
    #480.0; ADDR = 16'h20E9;
    #10.0; ADDR = 16'hA024;
    #410.0; ADDR = 16'hA025;
    #240.0; ADDR = 16'hA024;
    #10.0; ADDR = 16'hA026;
    #400.0; ADDR = 16'hA027;
    #410.0; ADDR = 16'hA028;
    #730.0; ADDR = 16'h9A00;
    #10.0; ADDR = 16'h1A97;
    #190.0; ADDR = 16'h1E97;
    #10.0; ADDR = 16'h1A97;
    #280.0; ADDR = 16'h2093;
    #10.0; ADDR = 16'hA029;
    #400.0; ADDR = 16'hA02B;
    #10.0; ADDR = 16'hA02A;
    #650.0; ADDR = 16'hA02F;
    #410.0; ADDR = 16'hA030;
    #410.0; ADDR = 16'hA031;
    #730.0; ADDR = 16'h2865;
    #10.0; ADDR = 16'h28E7;
    #320.0; ADDR = 16'hA032;
    #410.0; ADDR = 16'hA033;
    #410.0; ADDR = 16'hA034;
    #730.0; ADDR = 16'h1A10;
    #10.0; ADDR = 16'h1A9B;
    #480.0; ADDR = 16'h2033;
    #10.0; ADDR = 16'hA035;
    #400.0; ADDR = 16'hA037;
    #10.0; ADDR = 16'hA036;
    #490.0; ADDR = 16'hA037;
    #400.0; ADDR = 16'hA030;
    #10.0; ADDR = 16'hA038;
    #410.0; ADDR = 16'hA039;
    #720.0; ADDR = 16'h8039;
    #10.0; ADDR = 16'h1A9B;
    #570.0; ADDR = 16'hA03A;
    #410.0; ADDR = 16'hA03B;
    #410.0; ADDR = 16'hA03C;
    #730.0; ADDR = 16'h1A18;
    #10.0; ADDR = 16'h1A99;
    #570.0; ADDR = 16'h1A9A;
    #400.0; ADDR = 16'h209A;
    #10.0; ADDR = 16'hA03D;
    #400.0; ADDR = 16'hA03C;
    #10.0; ADDR = 16'hA03E;
    #410.0; ADDR = 16'hA03F;
    #160.0; ADDR = 16'h28E7;
    #570.0; ADDR = 16'h28E8;
    #400.0; ADDR = 16'h20E8;
    #10.0; ADDR = 16'hA03F;
    #410.0; ADDR = 16'hA040;
    #410.0; ADDR = 16'hA041;
    #730.0; ADDR = 16'h1A05;
    #10.0; ADDR = 16'h1A97;
    #480.0; ADDR = 16'h1A98;
    #410.0; ADDR = 16'h2042;
    #10.0; ADDR = 16'hA042;
    #400.0; ADDR = 16'hA043;
    #490.0; ADDR = 16'hA040;
    #10.0; ADDR = 16'hA044;
    #410.0; ADDR = 16'hA045;
    #640.0; ADDR = 16'h9845;
    #10.0; ADDR = 16'h1FED;
    #810.0; ADDR = 16'h1FEC;
    #410.0; ADDR = 16'h1FE8;
    #10.0; ADDR = 16'h1FEB;
    #230.0; ADDR = 16'h27EB;
    #10.0; ADDR = 16'hA046;
    #410.0; ADDR = 16'hA047;
    #650.0; ADDR = 16'h1FEC;
    #820.0; ADDR = 16'h1FED;
    #410.0; ADDR = 16'h1FEE;
    #320.0; ADDR = 16'h20EE;
    #10.0; ADDR = 16'hA048;
    #410.0; ADDR = 16'hA049;
    #400.0; ADDR = 16'hA048;
    #10.0; ADDR = 16'hA04A;
    #150.0; ADDR = 16'hA842;
    #10.0; ADDR = 16'h28E7;
    #570.0; ADDR = 16'h28E8;
    #400.0; ADDR = 16'h20E8;
    #10.0; ADDR = 16'hA04A;
    #410.0; ADDR = 16'hA04B;
    #400.0; ADDR = 16'hA048;
    #10.0; ADDR = 16'hA04C;
    #160.0; ADDR = 16'h020C;
    #900.0; ADDR = 16'h020D;
    #650.0; ADDR = 16'h200C;
    #10.0; ADDR = 16'hA04C;
    #400.0; ADDR = 16'hA04D;
    #160.0; ADDR = 16'h984D;
    #10.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h1FEF;
    #400.0; ADDR = 16'h1FF8;
    #10.0; ADDR = 16'h9FD8;
    #410.0; ADDR = 16'h9FD9;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDA;
    #730.0; ADDR = 16'h1A9C;
    #320.0; ADDR = 16'h1A98;
    #10.0; ADDR = 16'h9FDB;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDC;
    #410.0; ADDR = 16'h9FDD;
    #560.0; ADDR = 16'h8FDD;
    #10.0; ADDR = 16'h08F0;
    #890.0; ADDR = 16'h08D0;
    #10.0; ADDR = 16'h9FDE;
    #400.0; ADDR = 16'h9FDF;
    #660.0; ADDR = 16'h9FD6;
    #410.0; ADDR = 16'h9FD7;
    #650.0; ADDR = 16'h1FEF;
    #410.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h9FEF;
    #410.0; ADDR = 16'h9FF0;
    #410.0; ADDR = 16'h9FF1;
    #160.0; ADDR = 16'h1A9C;
    #570.0; ADDR = 16'h1A90;
    #10.0; ADDR = 16'h9FF1;
    #400.0; ADDR = 16'h9FF3;
    #10.0; ADDR = 16'h9FF2;
    #240.0; ADDR = 16'h9FF3;
    #410.0; ADDR = 16'h9FF4;
    #410.0; ADDR = 16'h9FF5;
    #160.0; ADDR = 16'h1A9C;
    #980.0; ADDR = 16'h9FF5;
    #410.0; ADDR = 16'h9FF6;
    #250.0; ADDR = 16'h9FF7;
    #400.0; ADDR = 16'h9FF8;
    #420.0; ADDR = 16'h9FF9;
    #730.0; ADDR = 16'h1A9F;
    #490.0; ADDR = 16'h1AA0;
    #410.0; ADDR = 16'h9FFA;
    #410.0; ADDR = 16'h9FFB;
    #400.0; ADDR = 16'h9FF8;
    #10.0; ADDR = 16'h9FFC;
    #730.0; ADDR = 16'h1AA1;
    #490.0; ADDR = 16'h9BBD;
    #10.0; ADDR = 16'h9FFD;
    #400.0; ADDR = 16'h9FFE;
    #410.0; ADDR = 16'h9FFF;
    #740.0; ADDR = 16'h1AA1;
    #480.0; ADDR = 16'h20A1;
    #10.0; ADDR = 16'hA000;
    #410.0; ADDR = 16'hA001;
    #490.0; ADDR = 16'hA002;
    #410.0; ADDR = 16'hA003;
    #650.0; ADDR = 16'hA015;
    #410.0; ADDR = 16'hA016;
    #490.0; ADDR = 16'hA017;
    #410.0; ADDR = 16'hA018;
    #410.0; ADDR = 16'hA019;
    #160.0; ADDR = 16'h1A9C;
    #650.0; ADDR = 16'h2018;
    #10.0; ADDR = 16'hA019;
    #400.0; ADDR = 16'hA01B;
    #10.0; ADDR = 16'hA01A;
    #400.0; ADDR = 16'hA01B;
    #730.0; ADDR = 16'h881B;
    #10.0; ADDR = 16'h1AA1;
    #480.0; ADDR = 16'h12A1;
    #10.0; ADDR = 16'hA01C;
    #410.0; ADDR = 16'hA01D;
    #240.0; ADDR = 16'hA01C;
    #10.0; ADDR = 16'hA01E;
    #400.0; ADDR = 16'hA01F;
    #410.0; ADDR = 16'hA020;
    #730.0; ADDR = 16'hA820;
    #10.0; ADDR = 16'h28F1;
    #320.0; ADDR = 16'h2021;
    #10.0; ADDR = 16'hA021;
    #400.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA022;
    #400.0; ADDR = 16'hA023;
    #730.0; ADDR = 16'hA823;
    #10.0; ADDR = 16'h28EF;
    #480.0; ADDR = 16'h20EF;
    #10.0; ADDR = 16'hA024;
    #410.0; ADDR = 16'hA025;
    #240.0; ADDR = 16'hA024;
    #10.0; ADDR = 16'hA026;
    #400.0; ADDR = 16'hA027;
    #410.0; ADDR = 16'hA028;
    #730.0; ADDR = 16'h9828;
    #10.0; ADDR = 16'h1A9D;
    #480.0; ADDR = 16'h209D;
    #10.0; ADDR = 16'hA029;
    #410.0; ADDR = 16'hA02A;
    #650.0; ADDR = 16'hA02F;
    #410.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA030;
    #400.0; ADDR = 16'hA031;
    #730.0; ADDR = 16'h2821;
    #10.0; ADDR = 16'h28ED;
    #320.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA032;
    #400.0; ADDR = 16'hA033;
    #410.0; ADDR = 16'hA034;
    #730.0; ADDR = 16'h9A20;
    #10.0; ADDR = 16'h1AA1;
    #480.0; ADDR = 16'h20A1;
    #10.0; ADDR = 16'hA035;
    #400.0; ADDR = 16'hA037;
    #10.0; ADDR = 16'hA036;
    #490.0; ADDR = 16'hA037;
    #400.0; ADDR = 16'hA038;
    #420.0; ADDR = 16'hA039;
    #730.0; ADDR = 16'h1AA1;
    #570.0; ADDR = 16'hA03A;
    #410.0; ADDR = 16'hA03B;
    #410.0; ADDR = 16'hA03C;
    #730.0; ADDR = 16'h1A1C;
    #10.0; ADDR = 16'h1A9F;
    #570.0; ADDR = 16'h1AA0;
    #400.0; ADDR = 16'h20A0;
    #10.0; ADDR = 16'hA03D;
    #400.0; ADDR = 16'hA03C;
    #10.0; ADDR = 16'hA03E;
    #410.0; ADDR = 16'hA03F;
    #150.0; ADDR = 16'hA83F;
    #10.0; ADDR = 16'h28ED;
    #570.0; ADDR = 16'h28EE;
    #400.0; ADDR = 16'h20EE;
    #10.0; ADDR = 16'hA03F;
    #410.0; ADDR = 16'hA040;
    #410.0; ADDR = 16'hA041;
    #730.0; ADDR = 16'h1A9D;
    #490.0; ADDR = 16'h1A9E;
    #120.0; ADDR = 16'h1E9E;
    #10.0; ADDR = 16'h1A9E;
    #280.0; ADDR = 16'hA042;
    #410.0; ADDR = 16'hA043;
    #490.0; ADDR = 16'hA044;
    #410.0; ADDR = 16'hA045;
    #650.0; ADDR = 16'h1F6D;
    #10.0; ADDR = 16'h1FED;
    #810.0; ADDR = 16'h1FEC;
    #410.0; ADDR = 16'h1FEB;
    #240.0; ADDR = 16'h2047;
    #10.0; ADDR = 16'hA046;
    #400.0; ADDR = 16'hA047;
    #650.0; ADDR = 16'h9847;
    #10.0; ADDR = 16'h1FEC;
    #820.0; ADDR = 16'h1FED;
    #400.0; ADDR = 16'h1FEE;
    #330.0; ADDR = 16'hA048;
    #410.0; ADDR = 16'hA049;
    #400.0; ADDR = 16'hA048;
    #10.0; ADDR = 16'hA04A;
    #160.0; ADDR = 16'h28EC;
    #10.0; ADDR = 16'h28ED;
    #560.0; ADDR = 16'h28EC;
    #10.0; ADDR = 16'h28EE;
    #400.0; ADDR = 16'hA04A;
    #410.0; ADDR = 16'hA04B;
    #410.0; ADDR = 16'hA04C;
    #160.0; ADDR = 16'h020E;
    #910.0; ADDR = 16'h020F;
    #640.0; ADDR = 16'h200C;
    #10.0; ADDR = 16'hA04C;
    #400.0; ADDR = 16'hA04D;
    #160.0; ADDR = 16'h804D;
    #10.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h1FEF;
    #400.0; ADDR = 16'h1FE8;
    #10.0; ADDR = 16'h9FD8;
    #410.0; ADDR = 16'h9FD9;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDA;
    #730.0; ADDR = 16'h1AA2;
    #320.0; ADDR = 16'h1A82;
    #10.0; ADDR = 16'h9FDB;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDC;
    #410.0; ADDR = 16'h9FDD;
    #560.0; ADDR = 16'h8FDD;
    #10.0; ADDR = 16'h08F0;
    #890.0; ADDR = 16'h08D0;
    #10.0; ADDR = 16'h9FDE;
    #410.0; ADDR = 16'h9FDF;
    #650.0; ADDR = 16'h9FD6;
    #410.0; ADDR = 16'h9FD7;
    #650.0; ADDR = 16'h1FCF;
    #10.0; ADDR = 16'h1FEF;
    #400.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h9FEF;
    #410.0; ADDR = 16'h9FF0;
    #410.0; ADDR = 16'h9FF1;
    #160.0; ADDR = 16'h1AA2;
    #570.0; ADDR = 16'h1AA0;
    #10.0; ADDR = 16'h9FF1;
    #400.0; ADDR = 16'h9FF3;
    #10.0; ADDR = 16'h9FF2;
    #240.0; ADDR = 16'h9FF3;
    #410.0; ADDR = 16'h9FF4;
    #410.0; ADDR = 16'h9FF5;
    #160.0; ADDR = 16'h1AA2;
    #980.0; ADDR = 16'h9FF4;
    #10.0; ADDR = 16'h9FF5;
    #400.0; ADDR = 16'h9FF6;
    #250.0; ADDR = 16'h9FF7;
    #400.0; ADDR = 16'h9FF8;
    #420.0; ADDR = 16'h9FF9;
    #730.0; ADDR = 16'h1AA5;
    #490.0; ADDR = 16'h1AA6;
    #400.0; ADDR = 16'h1AA2;
    #10.0; ADDR = 16'h9FFA;
    #410.0; ADDR = 16'h9FFB;
    #400.0; ADDR = 16'h9FF8;
    #10.0; ADDR = 16'h9FFC;
    #730.0; ADDR = 16'h1AA7;
    #490.0; ADDR = 16'h9FFD;
    #410.0; ADDR = 16'h9FFE;
    #410.0; ADDR = 16'h9FFF;
    #730.0; ADDR = 16'h1AA7;
    #490.0; ADDR = 16'h20A3;
    #10.0; ADDR = 16'hA000;
    #400.0; ADDR = 16'hA001;
    #490.0; ADDR = 16'hA000;
    #10.0; ADDR = 16'hA002;
    #410.0; ADDR = 16'hA003;
    #650.0; ADDR = 16'hA015;
    #400.0; ADDR = 16'hA014;
    #10.0; ADDR = 16'hA016;
    #490.0; ADDR = 16'hA017;
    #400.0; ADDR = 16'hA010;
    #10.0; ADDR = 16'hA018;
    #410.0; ADDR = 16'hA019;
    #150.0; ADDR = 16'h9819;
    #10.0; ADDR = 16'h1AA2;
    #650.0; ADDR = 16'hA019;
    #410.0; ADDR = 16'hA01A;
    #410.0; ADDR = 16'hA01B;
    #730.0; ADDR = 16'h1A03;
    #10.0; ADDR = 16'h1AA7;
    #190.0; ADDR = 16'h1EA7;
    #10.0; ADDR = 16'h1AA7;
    #280.0; ADDR = 16'h20AF;
    #10.0; ADDR = 16'hA01C;
    #400.0; ADDR = 16'hA01D;
    #250.0; ADDR = 16'hA01E;
    #410.0; ADDR = 16'hA01F;
    #400.0; ADDR = 16'hA017;
    #10.0; ADDR = 16'hA020;
    #730.0; ADDR = 16'h2820;
    #10.0; ADDR = 16'h28F7;
    #320.0; ADDR = 16'hA021;
    #410.0; ADDR = 16'hA022;
    #410.0; ADDR = 16'hA023;
    #730.0; ADDR = 16'h2821;
    #10.0; ADDR = 16'h28F5;
    #480.0; ADDR = 16'h2024;
    #10.0; ADDR = 16'hA024;
    #410.0; ADDR = 16'hA025;
    #240.0; ADDR = 16'hA026;
    #410.0; ADDR = 16'hA027;
    #400.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA028;
    #730.0; ADDR = 16'h1AA2;
    #10.0; ADDR = 16'h1AA3;
    #480.0; ADDR = 16'hA029;
    #410.0; ADDR = 16'hA02A;
    #660.0; ADDR = 16'hA02F;
    #400.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA030;
    #410.0; ADDR = 16'hA031;
    #730.0; ADDR = 16'h28F3;
    #320.0; ADDR = 16'h20F3;
    #10.0; ADDR = 16'hA032;
    #410.0; ADDR = 16'hA033;
    #400.0; ADDR = 16'hA030;
    #10.0; ADDR = 16'hA034;
    #730.0; ADDR = 16'h1AA7;
    #490.0; ADDR = 16'hA035;
    #410.0; ADDR = 16'hA036;
    #490.0; ADDR = 16'hA037;
    #410.0; ADDR = 16'hA038;
    #410.0; ADDR = 16'hA039;
    #730.0; ADDR = 16'h1AA7;
    #570.0; ADDR = 16'h2032;
    #10.0; ADDR = 16'hA03A;
    #400.0; ADDR = 16'hA03B;
    #410.0; ADDR = 16'hA03C;
    #730.0; ADDR = 16'h983C;
    #10.0; ADDR = 16'h1AA5;
    #570.0; ADDR = 16'h1AA6;
    #400.0; ADDR = 16'h02A6;
    #10.0; ADDR = 16'hA03D;
    #410.0; ADDR = 16'hA03E;
    #410.0; ADDR = 16'hA03F;
    #160.0; ADDR = 16'h28F3;
    #570.0; ADDR = 16'h28F0;
    #10.0; ADDR = 16'h28F4;
    #400.0; ADDR = 16'h2037;
    #10.0; ADDR = 16'hA03F;
    #400.0; ADDR = 16'hA000;
    #10.0; ADDR = 16'hA040;
    #400.0; ADDR = 16'hA041;
    #730.0; ADDR = 16'h1A01;
    #10.0; ADDR = 16'h1AA3;
    #490.0; ADDR = 16'h1AA4;
    #400.0; ADDR = 16'h20A4;
    #10.0; ADDR = 16'hA042;
    #400.0; ADDR = 16'hA043;
    #410.0; ADDR = 16'hB3C3;
    #10.0; ADDR = 16'hA043;
    #70.0; ADDR = 16'hA040;
    #10.0; ADDR = 16'hA044;
    #410.0; ADDR = 16'hA045;
    #640.0; ADDR = 16'h8045;
    #10.0; ADDR = 16'h1FED;
    #820.0; ADDR = 16'h1FEC;
    #400.0; ADDR = 16'h1FE8;
    #10.0; ADDR = 16'h1FEB;
    #240.0; ADDR = 16'hA046;
    #410.0; ADDR = 16'hA047;
    #650.0; ADDR = 16'h1B44;
    #10.0; ADDR = 16'h1FEC;
    #810.0; ADDR = 16'h1FED;
    #410.0; ADDR = 16'h1FEE;
    #320.0; ADDR = 16'h27EE;
    #10.0; ADDR = 16'hA048;
    #410.0; ADDR = 16'hA049;
    #410.0; ADDR = 16'hA04A;
    #160.0; ADDR = 16'h28F3;
    #570.0; ADDR = 16'h28F0;
    #10.0; ADDR = 16'h28F4;
    #400.0; ADDR = 16'hA042;
    #10.0; ADDR = 16'hA04A;
    #400.0; ADDR = 16'hA04B;
    #410.0; ADDR = 16'hA04C;
    #160.0; ADDR = 16'h0210;
    #910.0; ADDR = 16'h0211;
    #640.0; ADDR = 16'h2000;
    #10.0; ADDR = 16'hA04C;
    #400.0; ADDR = 16'hA04D;
    #160.0; ADDR = 16'h804D;
    #10.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h1FEF;
    #400.0; ADDR = 16'h1FE8;
    #10.0; ADDR = 16'h9FD8;
    #410.0; ADDR = 16'h9FD9;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDA;
    #730.0; ADDR = 16'h1AA8;
    #320.0; ADDR = 16'h1A88;
    #10.0; ADDR = 16'h9FDB;
    #400.0; ADDR = 16'h9FD8;
    #10.0; ADDR = 16'h9FDC;
    #410.0; ADDR = 16'h9FDD;
    #560.0; ADDR = 16'h8FFD;
    #10.0; ADDR = 16'h08F0;
    #890.0; ADDR = 16'h18D0;
    #10.0; ADDR = 16'h9FDE;
    #400.0; ADDR = 16'h9FDF;
    #660.0; ADDR = 16'h9FD6;
    #410.0; ADDR = 16'h9FD7;
    #650.0; ADDR = 16'h1FEF;
    #410.0; ADDR = 16'h1FEE;
    #410.0; ADDR = 16'h9FEF;
    #410.0; ADDR = 16'h9FF0;
    #410.0; ADDR = 16'h9FF1;
    #160.0; ADDR = 16'h1AA8;
    #570.0; ADDR = 16'h1AA0;
    #10.0; ADDR = 16'h9FF1;
    #400.0; ADDR = 16'h9FF2;
    #250.0; ADDR = 16'h9FF3;
    #410.0; ADDR = 16'h9FF4;
    #410.0; ADDR = 16'h9FF5;
    #160.0; ADDR = 16'h1AA8;
    #980.0; ADDR = 16'h9FF5;
    #410.0; ADDR = 16'h9FF6;
    #250.0; ADDR = 16'h9FF7;
    #400.0; ADDR = 16'h9FF8;
    #420.0; ADDR = 16'h9FF9;
    #730.0; ADDR = 16'h1AAB;
    #490.0; ADDR = 16'h1AAC;
    #410.0; ADDR = 16'h9FFA;
    #410.0; ADDR = 16'h9FFB;
    #410.0; ADDR = 16'h9FFC;
    #730.0; ADDR = 16'h1AAD;
    #500.0; ADDR = 16'h9FFD;
    #400.0; ADDR = 16'h9FFE;
    #410.0; ADDR = 16'h9FFF;
    #740.0; ADDR = 16'h1AAD;
    #480.0; ADDR = 16'h22AD;
    #10.0; ADDR = 16'hA000;
    #410.0; ADDR = 16'hA001;
    #490.0; ADDR = 16'hA002;
    #410.0; ADDR = 16'hA003;
    #650.0; ADDR = 16'hA015;
    #410.0; ADDR = 16'hA016;
    #490.0; ADDR = 16'hA017;
    #410.0; ADDR = 16'hA018;
    #410.0; ADDR = 16'hA019;
    #160.0; ADDR = 16'h1AA8;
    #650.0; ADDR = 16'h2009;
    #10.0; ADDR = 16'hA019;
    #400.0; ADDR = 16'hA01B;
    #10.0; ADDR = 16'hA01A;
    #400.0; ADDR = 16'hA01B;
    #730.0; ADDR = 16'h981B;
    #10.0; ADDR = 16'h1AAD;
    #200.0; ADDR = 16'h1EAD;
    #10.0; ADDR = 16'h1AAD;
    #270.0; ADDR = 16'h02AD;
    #10.0; ADDR = 16'hA01C;
    #410.0; ADDR = 16'hA01D;
    #240.0; ADDR = 16'hA01C;
    #10.0; ADDR = 16'hA01E;
    #410.0; ADDR = 16'hA01F;
    #400.0; ADDR = 16'hA020;
    #730.0; ADDR = 16'hA820;
    #10.0; ADDR = 16'h28FD;
    #320.0; ADDR = 16'h20E1;
    #10.0; ADDR = 16'hA021;
    #400.0; ADDR = 16'hA020;
    #10.0; ADDR = 16'hA022;
    #410.0; ADDR = 16'hA023;
    #730.0; ADDR = 16'h28FB;
    #480.0; ADDR = 16'h20FB;
    #10.0; ADDR = 16'hA024;
    #410.0; ADDR = 16'hA025;
    #240.0; ADDR = 16'hA024;
    #10.0; ADDR = 16'hA026;
    #410.0; ADDR = 16'hA027;
    #400.0; ADDR = 16'hA028;
    #730.0; ADDR = 16'h9828;
    #10.0; ADDR = 16'h1AA9;
    #480.0; ADDR = 16'h20A9;
    #10.0; ADDR = 16'hA029;
    #400.0; ADDR = 16'hA02B;
    #10.0; ADDR = 16'hA02A;
    #650.0; ADDR = 16'hA02F;
    #410.0; ADDR = 16'hA030;
    #410.0; ADDR = 16'hA031;
    #730.0; ADDR = 16'h2831;
    #10.0; ADDR = 16'h28F9;
    #320.0; ADDR = 16'hA032;
    #410.0; ADDR = 16'hA033;
    #410.0; ADDR = 16'hA034;
    #730.0; ADDR = 16'h1A24;
    #10.0; ADDR = 16'h1AAD;
    #480.0; ADDR = 16'h20A5;
    #10.0; ADDR = 16'hA035;
    #400.0; ADDR = 16'hA037;
    #10.0; ADDR = 16'hA036;
    #490.0; ADDR = 16'hA037;
    #400.0; ADDR = 16'hA030;
    #10.0; ADDR = 16'hA038;
    #410.0; ADDR = 16'hA039;
    #720.0; ADDR = 16'h8039;
    #10.0; ADDR = 16'h1AAD;
    #570.0; ADDR = 16'hA03A;
    #410.0; ADDR = 16'hA03B;
    #410.0; ADDR = 16'hA03C;
    #730.0; ADDR = 16'h1A28;
    #10.0; ADDR = 16'h1AAB;
    #570.0; ADDR = 16'h1AAC;
    #400.0; ADDR = 16'h20AC;
    #10.0; ADDR = 16'hA03D;
    #400.0; ADDR = 16'hA03C;
    #10.0; ADDR = 16'hA03E;
    #410.0; ADDR = 16'hA03F;
    #150.0; ADDR = 16'hA83F;
    #10.0; ADDR = 16'h28F9;
    #570.0; ADDR = 16'h28FA;
    #400.0; ADDR = 16'h20FA;
    #10.0; ADDR = 16'hA03F;
    #400.0; ADDR = 16'hA037;
    #10.0; ADDR = 16'hA040;
    #410.0; ADDR = 16'hA041;
    #730.0; ADDR = 16'h1AA9;
    #490.0; ADDR = 16'h1AAA;
    #120.0; ADDR = 16'h1EAA;
    #10.0; ADDR = 16'h1AAA;
    #280.0; ADDR = 16'hA042;
    #410.0; ADDR = 16'hA043;
    #490.0; ADDR = 16'hA044;
    #410.0; ADDR = 16'hA045;
    #650.0; ADDR = 16'h1F4D;
    #10.0; ADDR = 16'h1FED;
    #810.0; ADDR = 16'h1FEC;
    #410.0; ADDR = 16'h1FEB;
    #240.0; ADDR = 16'h20EB;
    #10.0; ADDR = 16'hA046;
    #400.0; ADDR = 16'hA047;
    #650.0; ADDR = 16'h8047;
    #10.0; ADDR = 16'h1FEC;
    #820.0; ADDR = 16'h1FED;
    #400.0; ADDR = 16'h1FEC;
    #10.0; ADDR = 16'h1FEE;
    #320.0; ADDR = 16'hA048;
    #410.0; ADDR = 16'hA049;
    #410.0; ADDR = 16'hA048;
    #10.0; ADDR = 16'hA04A;
    #150.0; ADDR = 16'h2848;
    #10.0; ADDR = 16'h28F9;
    #560.0; ADDR = 16'h28F8;
    #10.0; ADDR = 16'h28FA;
    #400.0; ADDR = 16'h204A;
    #10.0; ADDR = 16'hA04A;
    #410.0; ADDR = 16'hA04B;
    #400.0; ADDR = 16'hA048;
    #10.0; ADDR = 16'hA04C;
    #150.0; ADDR = 16'h0204;
    #10.0; ADDR = 16'h0212;
    #900.0; ADDR = 16'h0213;
    #640.0; ADDR = 16'h0013;
    #10.0; ADDR = 16'hA04C;
    #410.0; ADDR = 16'hA04D;
    #160.0; ADDR = 16'h1FEC;
    #10.0; ADDR = 16'h1FEE;
    #400.0; ADDR = 16'h1FEF;
    #410.0; ADDR = 16'h9FD8;
    #410.0; ADDR = 16'h9FD9;
    #410.0; ADDR = 16'h9FDA;
    #730.0; ADDR = 16'h1AAE;
    #330.0; ADDR = 16'h9F8B;
    #10.0; ADDR = 16'h9FDB;
    #400.0; ADDR = 16'h9FDC;
    #410.0; ADDR = 16'h9FDD;
    #570.0; ADDR = 16'h08F0;

end
initial
begin
    RWb = 1'b1;
    #9050.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #810.0; RWb = 1'b1;
    #6380.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5970.0; RWb = 1'b0;
    #1140.0; RWb = 1'b1;
    #5160.0; RWb = 1'b0;
    #400.0; RWb = 1'b1;
    #2130.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #3760.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #11290.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #16920.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #6370.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5970.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5150.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #2130.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #3760.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #11280.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #16930.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #810.0; RWb = 1'b1;
    #6380.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5970.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5150.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #2130.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #3760.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #11280.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #16930.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #1710.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #6380.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5960.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5150.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #2130.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #3760.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #11280.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #16920.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #6370.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5970.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5150.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #2130.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #3760.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #11280.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #16930.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #1710.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #6380.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;
    #5970.0; RWb = 1'b0;
    #1310.0; RWb = 1'b1;

end
initial
begin
    CRAMCS = 1'b1;
    #25770.0; CRAMCS = 1'b0;
    #370.0; CRAMCS = 1'b1;
    #290.0; CRAMCS = 1'b0;
    #370.0; CRAMCS = 1'b1;
    #58180.0; CRAMCS = 1'b0;
    #370.0; CRAMCS = 1'b1;
    #280.0; CRAMCS = 1'b0;
    #380.0; CRAMCS = 1'b1;
    #58180.0; CRAMCS = 1'b0;
    #370.0; CRAMCS = 1'b1;
    #280.0; CRAMCS = 1'b0;
    #380.0; CRAMCS = 1'b1;
    #58170.0; CRAMCS = 1'b0;
    #370.0; CRAMCS = 1'b1;
    #280.0; CRAMCS = 1'b0;
    #380.0; CRAMCS = 1'b1;
    #58170.0; CRAMCS = 1'b0;
    #370.0; CRAMCS = 1'b1;
    #280.0; CRAMCS = 1'b0;
    #380.0; CRAMCS = 1'b1;
    #58170.0; CRAMCS = 1'b0;
    #380.0; CRAMCS = 1'b1;
    #280.0; CRAMCS = 1'b0;
    #370.0; CRAMCS = 1'b1;

end
initial
begin
    DTAC2 = 1'b1;
    #10.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #690.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #360.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #440.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #850.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #690.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #370.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #850.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #690.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #850.0; DTAC2 = 1'b0;
    #90.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #370.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #440.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #690.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #370.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #850.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #690.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #440.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #370.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #440.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #690.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #360.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;

end
initial
begin
    AS = 1'b0;
    #200.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #570.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #580.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #320.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #410.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #250.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #90.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #420.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #320.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #580.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #570.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #250.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #90.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #570.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #580.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #250.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #420.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #570.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #580.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #320.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #250.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #420.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #580.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #570.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #250.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #730.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #80.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #330.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #500.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #160.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #570.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #580.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #170.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #320.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #410.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #330.0; AS = 1'b1;
    #490.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #80.0; AS = 1'b0;
    #570.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #250.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #740.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
    #90.0; AS = 1'b0;
    #320.0; AS = 1'b1;
end

endmodule